`timescale 1ns / 1ps

module and1(input logic a, b, output logic y);
        assign y = a & b;
        endmodule