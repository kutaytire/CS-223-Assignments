`timescale 1ns / 1ps


module notGate ( input logic a, output logic y);

assign y = ~a;
endmodule