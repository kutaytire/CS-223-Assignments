`timescale 1ns / 1ps

module FourToOneSim();

	logic d0,d1,d2,d3,s1,s2;
	logic y;

	FourToOneMuxStruc dut (d0,d1,d2,d3,s1,s2,y);

	initial begin

		d0 = 0; d1 = 0; d2 = 0; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d2 = 1; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d1 = 1; d2 = 0; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d2 = 1; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d0 = 1; d1 = 0; d2 = 0; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d2 = 1; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d1 = 1; d2 = 0; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d2 = 1; d3 = 0; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;
		d3 = 1; s1 = 0; s2 = 0; #10;
		s2 = 1; #10;
		s1 = 1; s2 = 0; #10;
		s2 = 1; #10;

	end
endmodule
