`timescale 1ns / 1ps

module xor1(input logic a, b, output logic y);
    assign y = a ^ b;
    endmodule