`timescale 1ns / 1ps

module inv ( input logic a, output logic y);

	assign y = ~a;
endmodule