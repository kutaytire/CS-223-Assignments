`timescale 1ns / 1ps

module or1(input logic a, b, output logic y);
            assign y = a | b;
            endmodule     