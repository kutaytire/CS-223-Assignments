`timescale 1ns / 1ps

module TestBenchComplex();

logic clk, reset, s1, s0, I0, I1, I2, I3, shr_in, shl_in;
logic  Q0, Q1, Q2, Q3;

MultiFunction dut (clk, reset, s1, s0, I0, I1, I2, I3, shr_in, shl_in, Q0, Q1, Q2, Q3);
   
   
   always 
    begin
    
     clk = 0; #5;
     clk = 1; #5;
    
    end
    initial begin 
    
    
        reset = 0;
        clk = 1;
        
        
        // s0 = 0 s1 = 0
        // shl_in = 0, shr_in = 0
        s0 = 0; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 0
        s0 = 0; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 0, shr_in = 1
        s0 = 0; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 1
        s0 = 0; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;        
        //s = 01
        // shl_in = 0, shr_in = 0
        s0 = 1; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 0
        s0 = 1; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 0, shr_in = 1
        s0 = 1; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 1
        s0 = 1; s1 = 0; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;   
        // s = 10 
        // shl_in = 0, shr_in = 0
        s0 = 0; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 0
        s0 = 0; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 0, shr_in = 1
        s0 = 0; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 1
        s0 = 0; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;   
        //s = 11 
        // shl_in = 0, shr_in = 0
        s0 = 1; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 0
        s0 = 1; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 0; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 0, shr_in = 1
        s0 = 1; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 0; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        //shl_in = 1, shr_in = 1
        s0 = 1; s1 = 1; I0 = 0; I1 = 0; I2 = 0; I3 = 0; shl_in = 1; shr_in = 1; #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I3 = 1; I2 = 0; I1 = 0; I0 = 0;                                             #10;
        I0 = 1;                                                                           #10;
        I1 = 1; I0 = 0;                                                                 #10;
        I0 = 1;                                                                           #10;
        I2 = 1; I1 = 0; I0 = 0;                                                       #10;
        I0 = 1;                                                                           #10;

	end
endmodule
